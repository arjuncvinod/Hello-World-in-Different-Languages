module hello;
  $display("Hello World");
endmodule
